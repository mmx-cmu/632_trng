`default_nettype none

module uart_ctl
  (input  logic clock, reset_n,
   output logic SCK, MOSI, SS);

    

endmodule : uart_ctl
