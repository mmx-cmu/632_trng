`default_nettype none

module uart_clk_gen
  #(parameter BASE_CLK = 25000000, BAUD=115200)
  (input  logic clk, reset_n,
   output logic clk2);

  logic [8:0] counter;

  always_ff @(posedge clk, negedge reset_n) begin
    if (~reset_n) begin
      counter <= 8'd433; //BASE_CLK/BAUD-1;
    end else begin
      counter <= counter - 1;
    end
  end

  assign clk2 = (counter == 8'b0);

endmodule : uart_clk_gen

module uart_ctl
  #(parameter BASE_CLK = 25000000, BAUD=115200)
  (input  logic       clk, reset_n,
   input  logic [7:0] bytes,
   input  logic       send,
   output logic       TX, done);

  logic uart_clk;
  uart_clk_gen #(.BASE_CLK(BASE_CLK), .BAUD(BAUD)) clk_gen(.clk, .reset_n, .clk2(uart_clk));

  /* shift register + counter for bits */
  logic counter_en, counter_clr;
  logic [3:0] counter;
  always_ff @(posedge uart_clk, posedge counter_clr) begin
    if (counter_clr) begin
      counter <= 4'd0;
    end else if (counter_en) begin
      counter <= counter + 1;
    end
  end

  // Automatically generated by ferris highroller on 2/21/2023, 2:56:11 PM
  enum logic [2:0] {
    WAIT_GO,
    SEND_START,
    SEND_BITS,
    SEND_STOP,
    DONE
  } cstate, nstate;

  always_comb begin
    nstate = cstate;
    done = 1'b0;
    TX = 1'b0;
    counter_en = 1'b0;
    counter_clr = 1'b0;

    case (cstate)
      WAIT_GO: begin
        TX = 1'b1;
        counter_clr = 1'b1;
        if (send) begin
          nstate = SEND_START;
        end
      end
      SEND_START: begin
        counter_en = 1'b1;
        TX = (counter < 4'd1);
        if (counter == 4'd2) begin
          nstate = SEND_BITS;
        end
      end
      SEND_BITS: begin
        TX = bytes[9 - counter];
        counter_en = 1'b1;
        if (counter == 4'd10) begin
          nstate = SEND_STOP;
          TX = 1'b1;
        end
      end
      SEND_STOP: begin
        TX = 1'b1;
        counter_en = 1'b1;
        if (counter == 4'd11) begin
          nstate = DONE;
        end
      end
      DONE: begin
        done = 1'b1;
        TX = 1'b1;
        counter_clr = 1'b1;
        if (~send) begin
          nstate = WAIT_GO;
        end
      end
    endcase
  end
  always_ff @(posedge clk, negedge reset_n) begin
    if (!reset_n) cstate <= WAIT_GO;
    else cstate <= nstate;
  end

endmodule : uart_ctl

`ifdef SIMULATION
module top();

  logic clk, reset_n, send, TX, done;
  logic [7:0] bytes;

  uart_ctl #(.BASE_CLK(500000)) dut(.*);

  initial begin
    reset_n = 1'b0;
    clk = 1'b0;
    #5 reset_n = 1'b1;
    forever #5 clk = ~clk;
  end

  initial begin
    bytes = 8'b1010_0110;
    send = 1'b0;
    @(posedge clk);
    @(posedge clk);
    send = 1'b1;
    @(posedge done);
    send = 1'b0;
    @(negedge done);
    bytes = 8'b1001_0101;
    send = 1'b1;
    @(posedge done);
    send = 1'b0;
    repeat (5000) @(posedge clk);
    bytes = 8'b1011_1101;
    send = 1'b1;
    @(posedge done);
    @(posedge clk);
    $finish();
  end

  initial begin
    #50000000 $display("timed out");
    $finish();
  end

endmodule : top
`endif
