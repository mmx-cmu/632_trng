`default_nettype none

//make sure we only send bits out at the agreed baudrate
//send a bit every 434 cycles (115200 bits/s)
module uart_clk_gen
  #(parameter BASE_CLK = 50000000, BAUD=115200)
  (input  logic clk, reset_n,
   output logic clk2);

  logic [15:0] counter;
  always_ff @(posedge clk, negedge reset_n) begin
    if (~reset_n) begin
      counter <= BASE_CLK/BAUD - 1;
    end else begin
      if (counter[15]) begin
        /* check if there is underflow */
        counter <= BASE_CLK/BAUD - 1;
      end else begin
        /* no underflow, keep going */
        counter <= counter - 1;
      end
    end
  end

  assign clk2 = (counter == 16'd0);

endmodule : uart_clk_gen

module uart_ctl
  #(parameter BASE_CLK = 50000000, BAUD=115200)
  (input  logic       clk, reset_n,
   input  logic [7:0] bits,
   input  logic       send,
   output logic       TX, done);

  logic uclk, uclk_rst;
  uart_clk_gen #(.BASE_CLK(BASE_CLK), .BAUD(BAUD)) clk_gen(.clk,
                                                           .reset_n(uclk_rst),
                                                           .clk2(uclk));

  // Automatically generated by ferris highroller on 2/21/2023, 9:54:11 PM
  enum logic [3:0] {
    WAIT_GO,
    SEND_START,
    SEND_BIT0,
    SEND_STOP,
    DONE,
    SEND_BIT1,
    SEND_BIT2,
    SEND_BIT3,
    SEND_BIT4,
    SEND_BIT5,
    SEND_BIT6,
    SEND_BIT7
  } cstate, nstate;
  
  always_comb begin
    nstate = cstate;
    uclk_rst = 1'b1;
    done = 1'b0;
    TX = 1'b0;
    
    case (cstate)
      WAIT_GO: begin
        TX = 1'b1;
        if (send) begin
          uclk_rst = 1'b0;
          nstate = SEND_START;
        end
      end
      SEND_START: begin
        if (uclk) begin
          nstate = SEND_BIT0;
        end
      end
      SEND_STOP: begin
        TX = 1'b1;
        if (uclk) begin
          nstate = DONE;
        end
      end
      DONE: begin
        done = 1'b1;
        TX = 1'b1;
        if (~send) begin
          nstate = WAIT_GO;
        end
      end
      SEND_BIT0: begin
        TX = bits[0];
        if (uclk) begin
          nstate = SEND_BIT1;
        end
      end
      SEND_BIT1: begin
        TX = bits[1];
        if (uclk) begin
          nstate = SEND_BIT2;
        end
      end
      SEND_BIT2: begin
        TX = bits[2];
        if (uclk) begin
          nstate = SEND_BIT3;
        end
      end
      SEND_BIT3: begin
        TX = bits[3];
        if (uclk) begin
          nstate = SEND_BIT4;
        end
      end
      SEND_BIT4: begin
        TX = bits[4];
        if (uclk) begin
          nstate = SEND_BIT5;
        end
      end
      SEND_BIT5: begin
        TX = bits[5];
        if (uclk) begin
          nstate = SEND_BIT6;
        end
      end
      SEND_BIT6: begin
        TX = bits[6];
        if (uclk) begin
          nstate = SEND_BIT7;
        end
      end
      SEND_BIT7: begin
        TX = bits[7];
        if (uclk) begin
          nstate = SEND_STOP;
        end
      end
    endcase
  end
  always_ff @(posedge clk, negedge reset_n) begin
    if (!reset_n) cstate <= WAIT_GO;
    else cstate <= nstate;
  end

endmodule : uart_ctl

`ifdef SIMULATION
module top();

  logic clk, reset_n, send, TX, done;
  logic [7:0] bits;

  uart_ctl dut(.*);

  initial begin
    reset_n = 1'b0;
    clk = 1'b0;
    #5 reset_n = 1'b1;
    forever #5 clk = ~clk;
  end

  initial begin
    bits = 8'b0001_0000;
    send = 1'b0;
    @(posedge clk);
    @(posedge clk);
    send = 1'b1;
    @(posedge done);
    send = 1'b0;
    @(negedge done);
    bits = 8'b1001_0101;
    send = 1'b1;
    @(posedge done);
    send = 1'b0;
    repeat (5000) @(posedge clk);
    bits = 8'b1011_1101;
    send = 1'b1;
    @(posedge done);
    @(posedge clk);
    $finish();
  end

  initial begin
    #50000000 $display("timed out");
    $finish();
  end

endmodule : top
`endif
